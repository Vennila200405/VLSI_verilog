module arithmetic_shift_right (
  input  wire signed [7:0] in,      
assign out = in >>> shift_amt;

endmodule
